module instruction_register(inst, );
	input [15:0] inst;
	
	
endmodule
