library verilog;
use verilog.vl_types.all;
entity testConroller is
end testConroller;
