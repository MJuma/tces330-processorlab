library verilog;
use verilog.vl_types.all;
entity test_program_counter is
end test_program_counter;
