library verilog;
use verilog.vl_types.all;
entity testProcessor is
end testProcessor;
