library verilog;
use verilog.vl_types.all;
entity test_Mux2_1 is
end test_Mux2_1;
