library verilog;
use verilog.vl_types.all;
entity testInstruction_register is
end testInstruction_register;
