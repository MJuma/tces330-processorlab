/*
This is just a test

*/
module LabB();


endmodule